library IEEE; 
use IEEE.STD_LOGIC_1164.all; 

entity ext16 is	--function extension
	port (a: in  STD_LOGIC_VECTOR (15 downto 0); 
		  y: out STD_LOGIC_VECTOR (31 downto 0)); 
end;

architecture behave of ext16 is 
begin 
	y <= a(15 downto 0) & x"0000"; 
end;